library verilog;
use verilog.vl_types.all;
entity test_johnson_counter is
end test_johnson_counter;
