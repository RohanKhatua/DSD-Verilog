library verilog;
use verilog.vl_types.all;
entity test_sipo is
end test_sipo;
