library verilog;
use verilog.vl_types.all;
entity test_jkff is
end test_jkff;
