library verilog;
use verilog.vl_types.all;
entity test_decade_counter is
end test_decade_counter;
