library verilog;
use verilog.vl_types.all;
entity test_add_sub is
end test_add_sub;
