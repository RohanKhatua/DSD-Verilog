library verilog;
use verilog.vl_types.all;
entity test_pipo is
end test_pipo;
