library verilog;
use verilog.vl_types.all;
entity test_ring_counter is
end test_ring_counter;
