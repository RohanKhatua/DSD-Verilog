library verilog;
use verilog.vl_types.all;
entity test_siso is
end test_siso;
