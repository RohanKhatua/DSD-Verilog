library verilog;
use verilog.vl_types.all;
entity test_mealy_fsm is
end test_mealy_fsm;
