library verilog;
use verilog.vl_types.all;
entity piso_test is
end piso_test;
